package fifo_shared_pkg;
    int NUM_TEST_CASES = 500;

    int error_count = 0;
    int correct_count = 0;
    bit test_finished = 0;

    event sample_event;
endpackage : fifo_shared_pkg