package fifo_transaction_pkg;

class fifo_transaction #(parameter FIFO_WIDTH = 16, FIFO_DEPTH = 8);
    rand bit rst_n;
    rand bit wr_en;
    rand bit rd_en;
    rand bit [FIFO_WIDTH-1:0] data_in;
    logic [FIFO_WIDTH-1:0] data_out;
    logic wr_ack;
    logic full;
    logic empty; 
    logic almostfull; 
    logic almostempty; 
    logic overflow;
    logic underflow;

    int RD_EN_ON_DIST, WR_EN_ON_DIST;

    function new (int rd_dist = 30, int wr_dist  = 70);
        this.RD_EN_ON_DIST = rd_dist;
        this.WR_EN_ON_DIST = wr_dist;
    endfunction

    constraint c_rst_n {
        rst_n dist {1 := 95, 0 := 5};
    }
    
    constraint c_wr_en {
        wr_en dist {1 := WR_EN_ON_DIST, 0 := (100 - WR_EN_ON_DIST)};
    }
    
    constraint c_rd_en {
        rd_en dist {1 := RD_EN_ON_DIST, 0 := (100 - RD_EN_ON_DIST)};
    }

    function string convert2string();
        return $sformatf("rst_n = %0b, wr_en = %0b, rd_en = %0b, data_in = 0x%0h, data_out = 0x%0h, wr_ack = %0b, full = %0b, empty = %0b, almostfull = %0b, almostempty = %0b, overflow = %0b, underflow = %0b", 
            rst_n, wr_en, rd_en, data_in, data_out, wr_ack, full, empty, almostfull, almostempty, overflow, underflow);
    endfunction
endclass : fifo_transaction

endpackage : fifo_transaction_pkg