import testing_pkg::*;

module ALU_tb;
    
endmodule